
/*
 * Transistor logic: output, input, control
 * PNP: drain, source, gate
 * NPN: source, drain, gate
 *
 * IHS <3
 */

module gate_xor (inp1, inp2, out);

    supply0 gnd;
    supply1 vdd;

    input  inp1;
    input  inp2;
    output out ;

    
    
endmodule


