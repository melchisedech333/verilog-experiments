
/*
 * Transistor logic: output, input, control
 * PNP: drain, source, gate
 * NPN: source, drain, gate
 *
 * IHS <3
 */

module half_adder (inp1, inp2, out, carry);

    supply0 gnd;
    supply1 vdd;

    input  inp1;
    input  inp2;
    output out;
    output carry;

    

endmodule


